`ifndef RAM_DEFINES
`define RAM_DEFINES

`define ADDR_WIDTH  9
`define DATA_WIDTH  32

`endif